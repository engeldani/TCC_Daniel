module tb_rodada;

endmodule
